* ECSE 330 SPICE PROJECT
* Christian Gallai - 260218797
* CKT Model w/ Ideal Op-Amp
* Analysis 2 - Frequency Response using a 1V AC input signal level

* Circuit Description

R1 1 2 8k
R2 2 3 8k
R3 3 4 10k
R4 2 7 10k
R5 5 6 10k
R6 6 7 10k
C1 2 3 9uF
C2 4 5 2uF
E1 3 0 0 2 1E6
E2 5 0 0 4 1E6
E3 7 0 0 6 1E6

Vi 1 0 AC 1V

* Analysis Request

.ac dec 5 10m 1k

*Output Request
.plot AC V(3)
.probe
.end